package alsu_test_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import alsu_env_pkt::*;  
  import alsu_config_pkg::*; 
  import alsu_reset_sequence_pkt::*; 
  import alsu_main_sequence_pkt::*; 

  class alsu_test extends uvm_test;
    `uvm_component_utils(alsu_test)

    alsu_env env;
    alsu_config alsu_cfg;
	virtual alu_if alsu_vif;
	alsu_reset_sequence reset_seq;
	alsu_main_sequence main_seq;

    function new(string name = "alsu_test", uvm_component parent = null);
      super.new(name, parent);
    endfunction

    function void build_phase(uvm_phase phase);
      super.build_phase(phase);
      env = alsu_env::type_id::create("env", this);
      alsu_cfg = alsu_config::type_id::create("alsu_cfg", this);
	  reset_seq = alsu_reset_sequence::type_id::create("reset_seq", this);
	  main_seq = alsu_main_sequence::type_id::create("main_seq", this);
      if (!uvm_config_db#(virtual alu_if)::get(this, "", "ALU_IF", alsu_cfg.alsu_vif))
        `uvm_fatal("build_phase", "Unable to get the virtual interface from uvm_config_db");
      uvm_config_db#(alsu_config)::set(this, "*", "CFG", alsu_cfg);
    endfunction

    task run_phase(uvm_phase phase);
      super.run_phase(phase);
      phase.raise_objection(this);
	  `uvm_info("run_phase","RESET ASSERTION.",UVM_LOW)
  reset_seq.start(env.agt.sqr);
	  `uvm_info("run_phase","RESET DEASSERTION.",UVM_LOW)
	  
	  `uvm_info("run_phase","STIMULUS START.",UVM_LOW)
      main_seq.start(env.agt.sqr);
      `uvm_info("run_phase","STIMULUS END.",UVM_LOW)

      phase.drop_objection(this);
    endtask

  endclass
endpackage


