
package alsu_env_pkt;
import uvm_pkg::*;
`include "uvm_macros.svh"

import alsu_agent_pkt::*;
import alsu_scoreboard_pkt::*;
import alsu_coverage_pkt::*;
import mysequencer_pkt::*;
class alsu_env extends uvm_env;
   `uvm_component_utils(alsu_env)
   
   alsu_agent agt;
   alsu_scoreboard sb;
   alsu_coverage cov;
   mysequencer seqr;
   function new(string name = "alsu_env", uvm_component parent = null);
      super.new(name, parent);
   endfunction
   
   function void build_phase(uvm_phase phase);
      super.build_phase(phase);
      agt = alsu_agent::type_id::create("agt", this);
      sb = alsu_scoreboard::type_id::create("sb", this);
      cov = alsu_coverage::type_id::create("cov", this);
       seqr = mysequencer::type_id::create("seqr", this);
   endfunction // build_phase
   
   function void connect_phase(uvm_phase phase);
      agt.agt_ap.connect(sb.sb_export);
      agt.agt_ap.connect(cov.cov_export);
   endfunction
endclass
endpackage